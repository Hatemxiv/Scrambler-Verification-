
package scr_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "scr_sequence_item.svh"
    `include "scr_sequence.svh"
    `include "scr_sequencer.svh"
    `include "scr_driver.svh"
    `include "scr_monitor.svh"
    `include "scr_agent.svh"
    `include "scr_scoreboard.svh"
    `include "scr_env.svh"
    `include "scr_test.svh"
    
endpackage: scr_pkg
